library verilog;
use verilog.vl_types.all;
entity DataPath_vlg_vec_tst is
end DataPath_vlg_vec_tst;
